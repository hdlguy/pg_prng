// This block implements LFSR polynomials from Xilinx document XAPP052.
module lfsr #(  
    parameter WIDTH = 16
) (  
    input   logic   [WIDTH-1:0]   datain,
    output  logic   [WIDTH-1:0]   dataout
);

    // this table is from Xilinx XAPP052
    const logic [3:64][63:0] coeff = '{
        64'h0000000000000006, // 3
        64'h000000000000000c, // 4
        64'h0000000000000014, // 5
        64'h0000000000000030, // 6
        64'h0000000000000060, // 7
        64'h00000000000000b8, // 8
        64'h0000000000000110, // 9
        64'h0000000000000240, // 10
        64'h0000000000000500, // 11
        64'h0000000000000829, // 12
        64'h000000000000100d, // 13
        64'h0000000000002015, // 14
        64'h0000000000006000, // 15
        64'h000000000000d008, // 16
        64'h0000000000012000, // 17
        64'h0000000000020400, // 18
        64'h0000000000040023, // 19
        64'h0000000000090000, // 20
        64'h0000000000140000, // 21
        64'h0000000000300000, // 22
        64'h0000000000420000, // 23
        64'h0000000000e10000, // 24
        64'h0000000001200000, // 25
        64'h0000000002000023, // 26
        64'h0000000004000013, // 27
        64'h0000000009000000, // 28
        64'h0000000014000000, // 29
        64'h0000000020000029, // 30
        64'h0000000048000000, // 31
        64'h0000000080200003, // 32
        64'h0000000100080000, // 33
        64'h0000000204000003, // 34
        64'h0000000500000000, // 35
        64'h0000000801000000, // 36
        64'h000000100000001f, // 37
        64'h0000002000000031, // 38
        64'h0000004400000000, // 39
        64'h000000a000140000, // 40
        64'h0000012000000000, // 41
        64'h00000300000c0000, // 42
        64'h0000063000000000, // 43
        64'h00000c0000030000, // 44
        64'h00001b0000000000, // 45
        64'h0000300003000000, // 46
        64'h0000420000000000, // 47
        64'h0000c00000180000, // 48
        64'h0001008000000000, // 49
        64'h0003000000c00000, // 50
        64'h0006000c00000000, // 51
        64'h0009000000000000, // 52
        64'h0018003000000000, // 53
        64'h0030000000030000, // 54
        64'h0040000040000000, // 55
        64'h00c0000600000000, // 56
        64'h0102000000000000, // 57
        64'h0200004000000000, // 58
        64'h0600003000000000, // 59
        64'h0c00000000000000, // 60
        64'h1800300000000000, // 61
        64'h3000000000000030, // 62
        64'h6000000000000000, // 63
        64'hd800000000000000  // 64
    };

    logic [WIDTH-1:0] xor_vec;
    assign xor_vec = (datain[0]) ? coeff[WIDTH][WIDTH-1:0] : 0;
    assign dataout = (datain>>1)^xor_vec;
    
endmodule: lfsr
                            

